magic
tech sky130A
magscale 1 2
timestamp 1715866809
<< viali >>
rect 248 7958 344 8024
rect 5630 7560 5732 7610
rect 5594 5904 5740 5958
<< metal1 >>
rect 132 14754 388 14998
rect 132 14694 376 14754
rect 183 14559 325 14694
rect 79 14417 325 14559
rect 79 13217 221 14417
rect -1780 8094 -1516 8106
rect -1780 8024 8256 8094
rect -1780 7958 248 8024
rect 344 7958 8256 8024
rect -1780 7894 8256 7958
rect -1780 7844 -1516 7894
rect 5078 7400 5310 7894
rect 5610 7610 5750 7894
rect 6182 7886 6229 7894
rect 5610 7560 5630 7610
rect 5732 7560 5750 7610
rect 5610 7546 5750 7560
rect 5642 7500 6150 7502
rect 5642 7466 6229 7500
rect 6182 7455 6229 7466
rect 5078 7234 5660 7400
rect 5920 7398 6084 7401
rect 5700 7395 6084 7398
rect 5700 7234 5920 7395
rect 5920 7228 6084 7234
rect 6182 7180 6228 7455
rect 6166 7177 6172 7180
rect 6093 7172 6172 7177
rect 5642 7136 6172 7172
rect 6093 7131 6172 7136
rect 6166 7128 6172 7131
rect 6224 7128 6230 7180
rect -1744 6762 -1480 6788
rect -1744 6570 8848 6762
rect -1744 6562 -1260 6570
rect -506 6562 -436 6570
rect -1744 6526 -1480 6562
rect 1119 6160 1294 6183
rect 1119 950 1294 5985
rect 5074 5760 5310 6570
rect 5571 6045 5757 6570
rect 6388 6052 6394 6260
rect 6602 6052 7442 6260
rect 5573 5958 5755 6045
rect 5573 5904 5594 5958
rect 5740 5904 5755 5958
rect 5573 5897 5755 5904
rect 6774 5858 6826 5864
rect 5630 5814 6774 5850
rect 5074 5596 5642 5760
rect 5850 5758 5928 5774
rect 5116 5590 5642 5596
rect 5684 5626 5928 5758
rect 6076 5626 6082 5774
rect 6172 5770 6208 5814
rect 6774 5800 6826 5806
rect 5684 5586 5918 5626
rect 6172 5542 6210 5770
rect 5628 5504 6210 5542
rect 7234 2520 7442 6052
rect 56 809 1294 950
rect 5284 2312 7442 2520
rect 56 778 1292 809
rect 1120 776 1292 778
rect 5284 -588 5492 2312
rect 5276 -796 5492 -588
<< via1 >>
rect 5920 7234 6084 7395
rect 6172 7128 6224 7180
rect 1119 5985 1294 6160
rect 6394 6052 6602 6260
rect 5928 5626 6076 5774
rect 6774 5806 6826 5858
<< metal2 >>
rect 1119 11109 1294 11118
rect 1119 6160 1294 10934
rect 5914 7234 5920 7395
rect 6084 7234 6090 7395
rect 5922 6926 6083 7234
rect 6172 7180 6224 7186
rect 6224 7167 6819 7168
rect 6903 7167 6912 7179
rect 6224 7131 6912 7167
rect 6172 7122 6224 7128
rect 6782 7130 6912 7131
rect 5928 6260 6076 6926
rect 6394 6260 6602 6266
rect 1113 5985 1119 6160
rect 1294 5985 1300 6160
rect 5920 6052 6394 6260
rect 5928 5774 6076 6052
rect 6394 6046 6602 6052
rect 6782 5858 6819 7130
rect 6903 7119 6912 7130
rect 6972 7119 6981 7179
rect 6768 5806 6774 5858
rect 6826 5806 6832 5858
rect 5928 5620 6076 5626
<< via2 >>
rect 1119 10934 1294 11109
rect 6912 7119 6972 7179
<< metal3 >>
rect 1114 11114 1299 11120
rect 1114 10934 1119 10939
rect 1294 10934 1299 10939
rect 1114 10929 1299 10934
rect 6907 7179 6977 7184
rect 7874 7179 7880 7181
rect 6907 7119 6912 7179
rect 6972 7119 7880 7179
rect 6907 7114 6977 7119
rect 7874 7117 7880 7119
rect 7944 7179 7950 7181
rect 7944 7119 7996 7179
rect 7944 7117 7950 7119
<< via3 >>
rect 1114 11109 1299 11114
rect 1114 10939 1119 11109
rect 1119 10939 1294 11109
rect 1294 10939 1299 11109
rect 7880 7117 7944 7181
<< metal4 >>
rect 1119 12768 5191 12943
rect 1119 11115 1294 12768
rect 1113 11114 1300 11115
rect 1113 10939 1114 11114
rect 1299 10939 1300 11114
rect 1113 10938 1300 10939
rect 7879 7181 7945 7182
rect 7879 7117 7880 7181
rect 7944 7179 7945 7181
rect 8766 7179 8826 9216
rect 7944 7119 8826 7179
rect 7944 7117 7945 7119
rect 7879 7116 7945 7117
use sky130_fd_pr__cap_mim_m3_1_BNHTNG  sky130_fd_pr__cap_mim_m3_1_BNHTNG_0
timestamp 1711880980
transform 1 0 6664 0 1 11124
box -2186 -2040 2186 2040
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1711880980
transform 1 0 5665 0 1 5676
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM2
timestamp 1711880980
transform 1 0 5679 0 1 7319
box -211 -319 211 319
use sky130_fd_pr__res_high_po_0p35_TTBX7G  XR1
timestamp 1711880980
transform 1 0 148 0 1 7129
box -201 -6582 201 6582
<< labels >>
flabel metal1 -1780 7844 -1516 8106 0 FreeSans 1600 0 0 0 vdd
port 4 nsew
flabel metal1 -1744 6526 -1480 6788 0 FreeSans 1600 0 0 0 vss
port 5 nsew
flabel metal1 5276 -796 5492 -588 0 FreeSans 1600 0 0 0 out
port 8 nsew
flabel metal1 132 14754 388 14998 0 FreeSans 1600 0 0 0 in
port 6 nsew
flabel metal2 1119 6160 1294 10934 0 FreeSans 1600 0 0 0 tocap
flabel metal3 6972 7119 7880 7179 0 FreeSans 1600 0 0 0 gate
<< end >>
